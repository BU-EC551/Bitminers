`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:31:50 03/03/2015 
// Design Name: 
// Module Name:    sync 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module sync(vga_h_sync, vga_v_sync, inDisplayArea, CounterX, CounterY,pixel_clk);
input pixel_clk;
output vga_h_sync, vga_v_sync;
output inDisplayArea;
output [9:0] CounterX;
output [8:0] CounterY;

//////////////////////////////////////////////////
<<<<<<< HEAD
initial 
begin
CounterX = 0;
CounterY= 0;
end

=======
>>>>>>> ca6f4445bd2340f9d05d89ab690fe74167c4cd9e
reg [9:0] CounterX;
reg [8:0] CounterY;
wire CounterXmaxed = (CounterX==10'h2FF);

always @(posedge pixel_clk)
if(CounterXmaxed)
	CounterX <= 0;
else
	CounterX <= CounterX + 1'b1;

always @(posedge pixel_clk)
if(CounterXmaxed) CounterY <= CounterY + 1'b1;

reg	vga_HS, vga_VS;
always @(posedge pixel_clk)
begin
	vga_HS <= (CounterX[9:4]==6'h2D); // change this value to move the display horizontally
	vga_VS <= (CounterY==500); // change this value to move the display vertically
end

reg inDisplayArea;
always @(posedge pixel_clk)
if(inDisplayArea==0)
	inDisplayArea <= (CounterXmaxed) && (CounterY<480);
else
	inDisplayArea <= !(CounterX==639);
	
assign vga_h_sync = ~vga_HS;
assign vga_v_sync = ~vga_VS;

endmodule
